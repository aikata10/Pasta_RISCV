`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/27/2020 06:50:26 PM
// Design Name: 
// Module Name: keccak_speed
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// Keccak HW architecture following the pseudocode algorithm specified in https://keccak.team/keccak_specs_summary.html

module keccak_speed(clk, rst, rounds_done,rateInBytes, delimitedSuffix, 
                inputLen_InBytes, outputLen_InBytes,
                keccak_is_ready_to_receive, din_64bit_raw, din_valid,
                keccak_squeeze_resume, dout_64bit, dout_valid, 
                absorb_done, squeeze_done);
input clk;
input rst,rounds_done;                      // Active high reset
input [7:0] rateInBytes;        // Note that maximum rateInBytes = 1344/8 = 168
input [7:0] delimitedSuffix;    // Keccak parameter    

input [15:0] inputLen_InBytes;  // Message length in bytes. If message is less than 64 bits, then the most significant bits are 0s.
input [15:0] outputLen_InBytes; // Length of output PRNG string in bytes.

output keccak_is_ready_to_receive;  // when this signal is high, that means Keccak is ready to absorb.
input [63:0] din_64bit_raw;
input din_valid;                    // This signal is provided by a data source to indicate that din_64bit_raw is valid

input keccak_squeeze_resume;     // This is used to 'resume' Keccak squeeze after a pause. Useful to generate PRNG in short chunks.
output [63:0] dout_64bit;        // 64-bit PRNG word output from Keccak state   
output dout_valid;               // This signal is used to write Keccak-squeeze output

output absorb_done; 
output squeeze_done;
//output done;                     // This signal goes 1 after requested Keccak (e.g., SHA, SHAKE) operation is completed


wire [63:0] din_64bit_processed;    // Properly padded message coming from keccak_absorb. It will be XORed with the State buffer.
wire din_wen;                       // This signal is generated by keccak_absorb to XOR din_64bit_processed with State.       
wire call_keccak_f1600_absorb;      // This is 1 to initiate F1600 on the state during Absorb. 
wire keccak_round_complete;         // Generated by Keccak-f1600 after it finishes a F1600.      
wire absorb_done;                   // Becomes 1 after the entire input message is absorbed.

wire [25*64-1:0] state_out;         // 25*64 bit state output from Keccak Buffer. It will be processed inside f1600 permutation.
wire [25*64-1:0] state_in;          // 25*64 bit new state value that will be written into the state bufer  
wire write_state_in;                // Write enable signal for writing the new state value into the state buffer. 

wire rst_f1600;

wire [4:0] state_reg_sel;           // This is used to select State[0]..to..State[rate] (at most). Note that only 64-bits are output every cycle.
wire we_output_buffer;       // Used to write keccak_state into keccak_output_buffer
wire shift_output_buffer;    // Used to shift the keccak_output_buffer in 64 bits such that one word is output
wire call_keccak_f1600_squeeze;     // This is 1 to initiate F1600 on the state during Squeeze
wire squeeze_done;             // Becomes 1 when the entire input is absorbed.

reg [2:0] FSM_state, FSM_nextstate;

reg rst_absorb, rst_state, rst_squeeze;
wire rst_rounds;
wire dout_valid_wire;

// Reset clears the state buffer.
// The first step is Keccak_absorb. This module is the FSM. It also does necessary padding to the message.
keccak_absorb Absorb(clk, rst_absorb, rateInBytes, inputLen_InBytes, delimitedSuffix,
                        din_64bit_raw, din_valid,
                        keccak_is_ready_to_receive, din_64bit_processed, din_wen, call_keccak_f1600_absorb,
                        keccak_round_complete, absorb_done);


keccak_state_buffer State(clk, rst_state, din_64bit_processed, din_wen, 
                            state_out, state_in, write_state_in, 
                            state_reg_sel, we_output_buffer, shift_output_buffer, dout_64bit);

assign rst_rounds = (rst_absorb==1'b0) ? ~call_keccak_f1600_absorb :
                    (rst_squeeze==1'b0) ? ~call_keccak_f1600_squeeze : 1'b1;
                    
keccak_f1600    Rounds(clk, rst_rounds, state_out, state_in, write_state_in, keccak_round_complete);


keccak_squeeze  Squeeze(clk, rounds_done,rst_squeeze, rateInBytes, outputLen_InBytes, keccak_squeeze_resume,
                        call_keccak_f1600_squeeze, keccak_round_complete, 
                        state_reg_sel, we_output_buffer, shift_output_buffer, dout_valid, squeeze_done);

//always @(posedge clk)
//    dout_valid <= dout_valid_wire;
    
always @(posedge clk)
begin
    if(rst)
        FSM_state <= 3'd0;
    else
        FSM_state <= FSM_nextstate;
end

always @(FSM_state)
begin
    case(FSM_state)
    3'd0: begin     // Reset state; Clear state buffer.
            rst_absorb<=1; rst_state<=1; rst_squeeze<=1;
         end

    3'd1: begin     // Absorb input
            rst_absorb<=0; rst_state<=0; rst_squeeze<=1;
         end

    3'd2: begin     // Squeeze
            rst_absorb<=1; rst_state<=0; rst_squeeze<=0;
         end

    3'd3: begin     // End state; Reset all.
            rst_absorb<=1; rst_state<=1; rst_squeeze<=1;
         end                  
    default: begin
            rst_absorb<=1; rst_state<=1; rst_squeeze<=1;
         end         
    endcase
end

always @(FSM_state or absorb_done or squeeze_done)
begin
    case(FSM_state)
    3'd0: FSM_nextstate <= 3'd1;

    3'd1: begin
            if(absorb_done)
                FSM_nextstate <= 3'd2;
            else
                FSM_nextstate <= 3'd1;
         end

    3'd2: begin
            if(squeeze_done)
                FSM_nextstate <= 3'd3;
            else
                FSM_nextstate <= 3'd2;
         end
         
    3'd3: FSM_nextstate <= 3'd3;
    default: FSM_nextstate <= 3'd0;    
    endcase
end

//assign done = (FSM_state==3'd3);

endmodule
